library verilog;
use verilog.vl_types.all;
entity processor_testbench is
end processor_testbench;
