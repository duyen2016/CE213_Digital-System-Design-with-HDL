library verilog;
use verilog.vl_types.all;
entity sram_tb is
end sram_tb;
